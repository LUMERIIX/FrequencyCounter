library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library work;
use work.zpupkg.all;
entity dualport_ram is

    generic(
        wordPower       : integer;
        maxAddrBitBRAM  : integer
    );
    port(
        clk             : in  std_logic;
        memAWriteEnable : in  std_logic;
        memAAddr        : in  std_logic_vector(maxAddrBitBRAM downto wordPower-3);
        memAWrite       : in  std_logic_vector(2**wordPower-1 downto 0);
        memARead        : out std_logic_vector(2**wordPower-1 downto 0);
        memBWriteEnable : in  std_logic;
        memBAddr        : in  std_logic_vector(maxAddrBitBRAM downto wordPower-3);
        memBWrite       : in  std_logic_vector(2**wordPower-1 downto 0);
        memBRead        : out std_logic_vector(2**wordPower-1 downto 0)
    );
end dualport_ram;

architecture dualport_ram_arch of dualport_ram is


    type ram_type is array(natural range 0 to ((2**(maxAddrBitBRAM+1))/4)-1) of std_logic_vector(2**wordPower-1 downto 0); 

    shared variable ram : ram_type :=
    (
             0 => x"0b0b0b9b",
             1 => x"e0040000",
             2 => x"00000000",
             3 => x"00000000",
             4 => x"00000000",
             5 => x"00000000",
             6 => x"00000000",
             7 => x"00000000",
             8 => x"0b0b0b89",
             9 => x"8f040000",
            10 => x"00000000",
            11 => x"00000000",
            12 => x"00000000",
            13 => x"00000000",
            14 => x"00000000",
            15 => x"00000000",
            16 => x"71fd0608",
            17 => x"72830609",
            18 => x"81058205",
            19 => x"832b2a83",
            20 => x"ffff0652",
            21 => x"04000000",
            22 => x"00000000",
            23 => x"00000000",
            24 => x"71fd0608",
            25 => x"83ffff73",
            26 => x"83060981",
            27 => x"05820583",
            28 => x"2b2b0906",
            29 => x"7383ffff",
            30 => x"0b0b0b0b",
            31 => x"83a70400",
            32 => x"72098105",
            33 => x"72057373",
            34 => x"09060906",
            35 => x"73097306",
            36 => x"070a8106",
            37 => x"53510400",
            38 => x"00000000",
            39 => x"00000000",
            40 => x"72722473",
            41 => x"732e0753",
            42 => x"51040000",
            43 => x"00000000",
            44 => x"00000000",
            45 => x"00000000",
            46 => x"00000000",
            47 => x"00000000",
            48 => x"71737109",
            49 => x"71068106",
            50 => x"30720a10",
            51 => x"0a720a10",
            52 => x"0a31050a",
            53 => x"81065151",
            54 => x"53510400",
            55 => x"00000000",
            56 => x"72722673",
            57 => x"732e0753",
            58 => x"51040000",
            59 => x"00000000",
            60 => x"00000000",
            61 => x"00000000",
            62 => x"00000000",
            63 => x"00000000",
            64 => x"00000000",
            65 => x"00000000",
            66 => x"00000000",
            67 => x"00000000",
            68 => x"00000000",
            69 => x"00000000",
            70 => x"00000000",
            71 => x"00000000",
            72 => x"0b0b0b88",
            73 => x"c3040000",
            74 => x"00000000",
            75 => x"00000000",
            76 => x"00000000",
            77 => x"00000000",
            78 => x"00000000",
            79 => x"00000000",
            80 => x"720a722b",
            81 => x"0a535104",
            82 => x"00000000",
            83 => x"00000000",
            84 => x"00000000",
            85 => x"00000000",
            86 => x"00000000",
            87 => x"00000000",
            88 => x"72729f06",
            89 => x"0981050b",
            90 => x"0b0b88a6",
            91 => x"05040000",
            92 => x"00000000",
            93 => x"00000000",
            94 => x"00000000",
            95 => x"00000000",
            96 => x"72722aff",
            97 => x"739f062a",
            98 => x"0974090a",
            99 => x"8106ff05",
           100 => x"06075351",
           101 => x"04000000",
           102 => x"00000000",
           103 => x"00000000",
           104 => x"71715351",
           105 => x"020d0406",
           106 => x"73830609",
           107 => x"81058205",
           108 => x"832b0b2b",
           109 => x"0772fc06",
           110 => x"0c515104",
           111 => x"00000000",
           112 => x"72098105",
           113 => x"72050970",
           114 => x"81050906",
           115 => x"0a810653",
           116 => x"51040000",
           117 => x"00000000",
           118 => x"00000000",
           119 => x"00000000",
           120 => x"72098105",
           121 => x"72050970",
           122 => x"81050906",
           123 => x"0a098106",
           124 => x"53510400",
           125 => x"00000000",
           126 => x"00000000",
           127 => x"00000000",
           128 => x"71098105",
           129 => x"52040000",
           130 => x"00000000",
           131 => x"00000000",
           132 => x"00000000",
           133 => x"00000000",
           134 => x"00000000",
           135 => x"00000000",
           136 => x"72720981",
           137 => x"05055351",
           138 => x"04000000",
           139 => x"00000000",
           140 => x"00000000",
           141 => x"00000000",
           142 => x"00000000",
           143 => x"00000000",
           144 => x"72097206",
           145 => x"73730906",
           146 => x"07535104",
           147 => x"00000000",
           148 => x"00000000",
           149 => x"00000000",
           150 => x"00000000",
           151 => x"00000000",
           152 => x"71fc0608",
           153 => x"72830609",
           154 => x"81058305",
           155 => x"1010102a",
           156 => x"81ff0652",
           157 => x"04000000",
           158 => x"00000000",
           159 => x"00000000",
           160 => x"71fc0608",
           161 => x"0b0b0b9d",
           162 => x"f0738306",
           163 => x"10100508",
           164 => x"060b0b0b",
           165 => x"88a90400",
           166 => x"00000000",
           167 => x"00000000",
           168 => x"0b0b0b88",
           169 => x"f7040000",
           170 => x"00000000",
           171 => x"00000000",
           172 => x"00000000",
           173 => x"00000000",
           174 => x"00000000",
           175 => x"00000000",
           176 => x"0b0b0b88",
           177 => x"df040000",
           178 => x"00000000",
           179 => x"00000000",
           180 => x"00000000",
           181 => x"00000000",
           182 => x"00000000",
           183 => x"00000000",
           184 => x"72097081",
           185 => x"0509060a",
           186 => x"8106ff05",
           187 => x"70547106",
           188 => x"73097274",
           189 => x"05ff0506",
           190 => x"07515151",
           191 => x"04000000",
           192 => x"72097081",
           193 => x"0509060a",
           194 => x"098106ff",
           195 => x"05705471",
           196 => x"06730972",
           197 => x"7405ff05",
           198 => x"06075151",
           199 => x"51040000",
           200 => x"05ff0504",
           201 => x"00000000",
           202 => x"00000000",
           203 => x"00000000",
           204 => x"00000000",
           205 => x"00000000",
           206 => x"00000000",
           207 => x"00000000",
           208 => x"810b0b0b",
           209 => x"0b9e940c",
           210 => x"51040000",
           211 => x"00000000",
           212 => x"00000000",
           213 => x"00000000",
           214 => x"00000000",
           215 => x"00000000",
           216 => x"71810552",
           217 => x"04000000",
           218 => x"00000000",
           219 => x"00000000",
           220 => x"00000000",
           221 => x"00000000",
           222 => x"00000000",
           223 => x"00000000",
           224 => x"00000000",
           225 => x"00000000",
           226 => x"00000000",
           227 => x"00000000",
           228 => x"00000000",
           229 => x"00000000",
           230 => x"00000000",
           231 => x"00000000",
           232 => x"02840572",
           233 => x"10100552",
           234 => x"04000000",
           235 => x"00000000",
           236 => x"00000000",
           237 => x"00000000",
           238 => x"00000000",
           239 => x"00000000",
           240 => x"00000000",
           241 => x"00000000",
           242 => x"00000000",
           243 => x"00000000",
           244 => x"00000000",
           245 => x"00000000",
           246 => x"00000000",
           247 => x"00000000",
           248 => x"717105ff",
           249 => x"05715351",
           250 => x"020d0400",
           251 => x"00000000",
           252 => x"00000000",
           253 => x"00000000",
           254 => x"00000000",
           255 => x"00000000",
           256 => x"82b03f95",
           257 => x"c03f0410",
           258 => x"10101010",
           259 => x"10101010",
           260 => x"10101010",
           261 => x"10101010",
           262 => x"10101010",
           263 => x"10101010",
           264 => x"10101010",
           265 => x"10105351",
           266 => x"047381ff",
           267 => x"06738306",
           268 => x"09810583",
           269 => x"05101010",
           270 => x"2b0772fc",
           271 => x"060c5151",
           272 => x"043c0472",
           273 => x"72807281",
           274 => x"06ff0509",
           275 => x"72060571",
           276 => x"1052720a",
           277 => x"100a5372",
           278 => x"ed385151",
           279 => x"53510480",
           280 => x"08840888",
           281 => x"08757599",
           282 => x"962d5050",
           283 => x"80085688",
           284 => x"0c840c80",
           285 => x"0c510480",
           286 => x"08840888",
           287 => x"08757597",
           288 => x"e42d5050",
           289 => x"80085688",
           290 => x"0c840c80",
           291 => x"0c510480",
           292 => x"08840888",
           293 => x"089ca02d",
           294 => x"880c840c",
           295 => x"800c049e",
           296 => x"9408802e",
           297 => x"a1389e98",
           298 => x"08822eb9",
           299 => x"38838080",
           300 => x"0b0b0b0b",
           301 => x"a6c40c82",
           302 => x"a0800ba6",
           303 => x"c80c8290",
           304 => x"800ba6cc",
           305 => x"0c04f880",
           306 => x"8080a40b",
           307 => x"0b0b0ba6",
           308 => x"c40cf880",
           309 => x"8082800b",
           310 => x"a6c80cf8",
           311 => x"80808480",
           312 => x"0ba6cc0c",
           313 => x"0480c0a8",
           314 => x"808c0b0b",
           315 => x"0b0ba6c4",
           316 => x"0c80c0a8",
           317 => x"80940ba6",
           318 => x"c80c9e80",
           319 => x"0ba6cc0c",
           320 => x"04ff3d0d",
           321 => x"a6d03351",
           322 => x"70a3389e",
           323 => x"a0087008",
           324 => x"52527080",
           325 => x"2e923884",
           326 => x"129ea00c",
           327 => x"702d9ea0",
           328 => x"08700852",
           329 => x"5270f038",
           330 => x"810ba6d0",
           331 => x"34833d0d",
           332 => x"0404803d",
           333 => x"0d0b0b0b",
           334 => x"a6c00880",
           335 => x"2e8e380b",
           336 => x"0b0b0b80",
           337 => x"0b802e09",
           338 => x"81068538",
           339 => x"823d0d04",
           340 => x"0b0b0ba6",
           341 => x"c0510b0b",
           342 => x"0bf5a53f",
           343 => x"823d0d04",
           344 => x"048c0802",
           345 => x"8c0cfc3d",
           346 => x"0d800b8c",
           347 => x"08fc050c",
           348 => x"800b8c08",
           349 => x"f8050c8c",
           350 => x"08fc0508",
           351 => x"8c08f405",
           352 => x"0c8c08f4",
           353 => x"0508812e",
           354 => x"b8388c08",
           355 => x"f4050881",
           356 => x"248c388c",
           357 => x"08f40508",
           358 => x"802e9938",
           359 => x"da398c08",
           360 => x"f4050882",
           361 => x"2e818738",
           362 => x"8c08f405",
           363 => x"08842e82",
           364 => x"e438c439",
           365 => x"84833f81",
           366 => x"0b8c08fc",
           367 => x"050cffb7",
           368 => x"399efc08",
           369 => x"70087087",
           370 => x"2a708106",
           371 => x"7081ff06",
           372 => x"51515151",
           373 => x"5170802e",
           374 => x"80ca389e",
           375 => x"c8089efc",
           376 => x"08700870",
           377 => x"83067074",
           378 => x"0c9ecc08",
           379 => x"9efc0870",
           380 => x"08708c06",
           381 => x"70822a70",
           382 => x"750c9ec0",
           383 => x"089efc08",
           384 => x"7008720c",
           385 => x"9ed00851",
           386 => x"52555151",
           387 => x"51525451",
           388 => x"51525280",
           389 => x"710c820b",
           390 => x"8c08fc05",
           391 => x"0c9ed408",
           392 => x"5181710c",
           393 => x"9efc0870",
           394 => x"085151fe",
           395 => x"ca399ed8",
           396 => x"08700870",
           397 => x"81067081",
           398 => x"ff065151",
           399 => x"51517080",
           400 => x"2efeb438",
           401 => x"9ed40851",
           402 => x"80710c9e",
           403 => x"ec087008",
           404 => x"70982b70",
           405 => x"81ff0a06",
           406 => x"a6f40c9e",
           407 => x"f0087008",
           408 => x"70902b70",
           409 => x"87fc8080",
           410 => x"0670a6f4",
           411 => x"0807a6f4",
           412 => x"0c9ef408",
           413 => x"70087088",
           414 => x"2b7083fe",
           415 => x"800670a6",
           416 => x"f40807a6",
           417 => x"f40c9ef8",
           418 => x"08700870",
           419 => x"81ff0670",
           420 => x"a6f40807",
           421 => x"a6f40c9e",
           422 => x"dc087008",
           423 => x"70982b70",
           424 => x"81ff0a06",
           425 => x"a6f80c9e",
           426 => x"e0087008",
           427 => x"70902b70",
           428 => x"87fc8080",
           429 => x"0670a6f8",
           430 => x"0807a6f8",
           431 => x"0c9ee408",
           432 => x"70087088",
           433 => x"2b7083fe",
           434 => x"800670a6",
           435 => x"f80807a6",
           436 => x"f80c9ee8",
           437 => x"08700870",
           438 => x"81ff0670",
           439 => x"a6f80807",
           440 => x"a6f80c51",
           441 => x"51515151",
           442 => x"51515151",
           443 => x"51515151",
           444 => x"51515151",
           445 => x"51515151",
           446 => x"51515151",
           447 => x"51515184",
           448 => x"0b8c08fc",
           449 => x"050c800b",
           450 => x"9f940c9e",
           451 => x"d0085181",
           452 => x"710cfce3",
           453 => x"399f8408",
           454 => x"70087081",
           455 => x"32708106",
           456 => x"7081ff06",
           457 => x"51515151",
           458 => x"5170802e",
           459 => x"fcc9389e",
           460 => x"d4085180",
           461 => x"710c9f94",
           462 => x"088738a6",
           463 => x"f4089f98",
           464 => x"0c9f9408",
           465 => x"842e0981",
           466 => x"068738a6",
           467 => x"f8089f98",
           468 => x"0c9f9408",
           469 => x"882e0981",
           470 => x"0696389f",
           471 => x"88085180",
           472 => x"710c9f80",
           473 => x"08518071",
           474 => x"0c810b8c",
           475 => x"08fc050c",
           476 => x"9efc0870",
           477 => x"087080f0",
           478 => x"0670842a",
           479 => x"51515151",
           480 => x"709f9408",
           481 => x"2e098106",
           482 => x"fbed389f",
           483 => x"80089f98",
           484 => x"08982a70",
           485 => x"720c9f88",
           486 => x"08515252",
           487 => x"81710c9f",
           488 => x"88085180",
           489 => x"710c9f98",
           490 => x"08882b9f",
           491 => x"980c9f94",
           492 => x"0881059f",
           493 => x"940cfbbf",
           494 => x"398c0802",
           495 => x"8c0cff3d",
           496 => x"0d9ea808",
           497 => x"5280720c",
           498 => x"9ea40852",
           499 => x"93720c9e",
           500 => x"ac085281",
           501 => x"80720c9e",
           502 => x"b0085280",
           503 => x"720c800b",
           504 => x"9f8c0c90",
           505 => x"80518a3f",
           506 => x"71800c83",
           507 => x"3d0d8c0c",
           508 => x"048c0802",
           509 => x"8c0cfe3d",
           510 => x"0d9ec008",
           511 => x"9ebc0870",
           512 => x"08720c52",
           513 => x"52800b8c",
           514 => x"08fc050c",
           515 => x"9f8c0851",
           516 => x"70832682",
           517 => x"da389f8c",
           518 => x"08517080",
           519 => x"c7389eb8",
           520 => x"08518190",
           521 => x"710c9eb0",
           522 => x"085181c8",
           523 => x"710c9ebc",
           524 => x"08700870",
           525 => x"812a7081",
           526 => x"067081ff",
           527 => x"06515151",
           528 => x"51517080",
           529 => x"2e8f388c",
           530 => x"08fc0508",
           531 => x"81058c08",
           532 => x"fc050cda",
           533 => x"39810b9f",
           534 => x"8c0c9ec4",
           535 => x"08518171",
           536 => x"0c81fd39",
           537 => x"9f8c0851",
           538 => x"70812e09",
           539 => x"8106bf38",
           540 => x"9eb00851",
           541 => x"80e0710c",
           542 => x"9eb80851",
           543 => x"90710c9e",
           544 => x"bc087008",
           545 => x"70812a70",
           546 => x"81067081",
           547 => x"ff065151",
           548 => x"51515170",
           549 => x"802e8f38",
           550 => x"8c08fc05",
           551 => x"0881058c",
           552 => x"08fc050c",
           553 => x"da39820b",
           554 => x"9f8c0c81",
           555 => x"b3399f8c",
           556 => x"08517082",
           557 => x"2e098106",
           558 => x"80c6389e",
           559 => x"b0088c08",
           560 => x"88050884",
           561 => x"2a70720c",
           562 => x"9eb80852",
           563 => x"53519071",
           564 => x"0c9ebc08",
           565 => x"70087081",
           566 => x"2a708106",
           567 => x"7081ff06",
           568 => x"51515151",
           569 => x"5170802e",
           570 => x"8f388c08",
           571 => x"fc050881",
           572 => x"058c08fc",
           573 => x"050cda39",
           574 => x"830b9f8c",
           575 => x"0c80e139",
           576 => x"9f8c0851",
           577 => x"70832e09",
           578 => x"810680d4",
           579 => x"389eb008",
           580 => x"8c088805",
           581 => x"088f0670",
           582 => x"842b7073",
           583 => x"0c9eb808",
           584 => x"51515252",
           585 => x"80d0710c",
           586 => x"9ebc0870",
           587 => x"0870812a",
           588 => x"70813270",
           589 => x"81067081",
           590 => x"ff065151",
           591 => x"51515151",
           592 => x"70802e8f",
           593 => x"388c08fc",
           594 => x"05088105",
           595 => x"8c08fc05",
           596 => x"0cd63984",
           597 => x"0b9f8c0c",
           598 => x"9eb80851",
           599 => x"80c0710c",
           600 => x"9ec0089e",
           601 => x"bc087008",
           602 => x"720c5252",
           603 => x"fd9e3980",
           604 => x"0b9f8c0c",
           605 => x"70800c84",
           606 => x"3d0d8c0c",
           607 => x"048c0802",
           608 => x"8c0cff3d",
           609 => x"0d800b8c",
           610 => x"08fc050c",
           611 => x"9ebc0870",
           612 => x"0870872a",
           613 => x"70813270",
           614 => x"81067081",
           615 => x"ff065151",
           616 => x"51515151",
           617 => x"70802eb8",
           618 => x"38a6e808",
           619 => x"5170b138",
           620 => x"9eb80851",
           621 => x"81a0710c",
           622 => x"9eb00851",
           623 => x"81c1710c",
           624 => x"9ebc0870",
           625 => x"0870812a",
           626 => x"70810670",
           627 => x"81ff0651",
           628 => x"51515151",
           629 => x"70802e83",
           630 => x"38e63981",
           631 => x"0ba6e80c",
           632 => x"9ebc0870",
           633 => x"0870872a",
           634 => x"70813270",
           635 => x"81067081",
           636 => x"ff065151",
           637 => x"51515151",
           638 => x"70802ebd",
           639 => x"38a6e808",
           640 => x"5170812e",
           641 => x"098106b1",
           642 => x"389eb808",
           643 => x"51a0710c",
           644 => x"9eb40870",
           645 => x"08a6dc0c",
           646 => x"519ebc08",
           647 => x"70087081",
           648 => x"2a708106",
           649 => x"7081ff06",
           650 => x"51515151",
           651 => x"5170802e",
           652 => x"8338e639",
           653 => x"820ba6e8",
           654 => x"0c9ebc08",
           655 => x"70087087",
           656 => x"2a708132",
           657 => x"70810670",
           658 => x"81ff0651",
           659 => x"51515151",
           660 => x"5170802e",
           661 => x"bd38a6e8",
           662 => x"08517082",
           663 => x"2e098106",
           664 => x"b1389eb8",
           665 => x"0851a071",
           666 => x"0c9eb408",
           667 => x"7008a6d4",
           668 => x"0c519ebc",
           669 => x"08700870",
           670 => x"812a7081",
           671 => x"067081ff",
           672 => x"06515151",
           673 => x"51517080",
           674 => x"2e8338e6",
           675 => x"39830ba6",
           676 => x"e80c9ebc",
           677 => x"08700870",
           678 => x"872a7081",
           679 => x"32708106",
           680 => x"7081ff06",
           681 => x"51515151",
           682 => x"51517080",
           683 => x"2ebd38a6",
           684 => x"e8085170",
           685 => x"832e0981",
           686 => x"06b1389e",
           687 => x"b80851a0",
           688 => x"710c9eb4",
           689 => x"087008a6",
           690 => x"d80c519e",
           691 => x"bc087008",
           692 => x"70812a70",
           693 => x"81067081",
           694 => x"ff065151",
           695 => x"51515170",
           696 => x"802e8338",
           697 => x"e639840b",
           698 => x"a6e80c9e",
           699 => x"bc087008",
           700 => x"70872a70",
           701 => x"81327081",
           702 => x"067081ff",
           703 => x"06515151",
           704 => x"51515170",
           705 => x"802ebd38",
           706 => x"a6e80851",
           707 => x"70842e09",
           708 => x"8106b138",
           709 => x"9eb80851",
           710 => x"a0710c9e",
           711 => x"b4087008",
           712 => x"a6e40c51",
           713 => x"9ebc0870",
           714 => x"0870812a",
           715 => x"70810670",
           716 => x"81ff0651",
           717 => x"51515151",
           718 => x"70802e83",
           719 => x"38e63985",
           720 => x"0ba6e80c",
           721 => x"9ebc0870",
           722 => x"0870872a",
           723 => x"70813270",
           724 => x"81067081",
           725 => x"ff065151",
           726 => x"51515151",
           727 => x"70802e80",
           728 => x"c538a6e8",
           729 => x"08517085",
           730 => x"2e098106",
           731 => x"b9389eb8",
           732 => x"0851a071",
           733 => x"0c9eb408",
           734 => x"7008a6e0",
           735 => x"0c519ebc",
           736 => x"08700870",
           737 => x"812a7081",
           738 => x"067081ff",
           739 => x"06515151",
           740 => x"51517080",
           741 => x"2e8338e6",
           742 => x"39800ba6",
           743 => x"e80c9eb8",
           744 => x"085180c0",
           745 => x"710ca6e8",
           746 => x"08517080",
           747 => x"2ead389e",
           748 => x"bc087008",
           749 => x"70862a70",
           750 => x"81327081",
           751 => x"067081ff",
           752 => x"06515151",
           753 => x"51515170",
           754 => x"802e9038",
           755 => x"9eb80851",
           756 => x"80c0710c",
           757 => x"9eb00851",
           758 => x"80710c70",
           759 => x"800c833d",
           760 => x"0d8c0c04",
           761 => x"8c08028c",
           762 => x"0cf93d0d",
           763 => x"800b8c08",
           764 => x"fc050c8c",
           765 => x"08880508",
           766 => x"8025ab38",
           767 => x"8c088805",
           768 => x"08308c08",
           769 => x"88050c80",
           770 => x"0b8c08f4",
           771 => x"050c8c08",
           772 => x"fc050888",
           773 => x"38810b8c",
           774 => x"08f4050c",
           775 => x"8c08f405",
           776 => x"088c08fc",
           777 => x"050c8c08",
           778 => x"8c050880",
           779 => x"25ab388c",
           780 => x"088c0508",
           781 => x"308c088c",
           782 => x"050c800b",
           783 => x"8c08f005",
           784 => x"0c8c08fc",
           785 => x"05088838",
           786 => x"810b8c08",
           787 => x"f0050c8c",
           788 => x"08f00508",
           789 => x"8c08fc05",
           790 => x"0c80538c",
           791 => x"088c0508",
           792 => x"528c0888",
           793 => x"05085181",
           794 => x"a73f8008",
           795 => x"708c08f8",
           796 => x"050c548c",
           797 => x"08fc0508",
           798 => x"802e8c38",
           799 => x"8c08f805",
           800 => x"08308c08",
           801 => x"f8050c8c",
           802 => x"08f80508",
           803 => x"70800c54",
           804 => x"893d0d8c",
           805 => x"0c048c08",
           806 => x"028c0cfb",
           807 => x"3d0d800b",
           808 => x"8c08fc05",
           809 => x"0c8c0888",
           810 => x"05088025",
           811 => x"93388c08",
           812 => x"88050830",
           813 => x"8c088805",
           814 => x"0c810b8c",
           815 => x"08fc050c",
           816 => x"8c088c05",
           817 => x"0880258c",
           818 => x"388c088c",
           819 => x"0508308c",
           820 => x"088c050c",
           821 => x"81538c08",
           822 => x"8c050852",
           823 => x"8c088805",
           824 => x"0851ad3f",
           825 => x"8008708c",
           826 => x"08f8050c",
           827 => x"548c08fc",
           828 => x"0508802e",
           829 => x"8c388c08",
           830 => x"f8050830",
           831 => x"8c08f805",
           832 => x"0c8c08f8",
           833 => x"05087080",
           834 => x"0c54873d",
           835 => x"0d8c0c04",
           836 => x"8c08028c",
           837 => x"0cfd3d0d",
           838 => x"810b8c08",
           839 => x"fc050c80",
           840 => x"0b8c08f8",
           841 => x"050c8c08",
           842 => x"8c05088c",
           843 => x"08880508",
           844 => x"27ac388c",
           845 => x"08fc0508",
           846 => x"802ea338",
           847 => x"800b8c08",
           848 => x"8c050824",
           849 => x"99388c08",
           850 => x"8c050810",
           851 => x"8c088c05",
           852 => x"0c8c08fc",
           853 => x"0508108c",
           854 => x"08fc050c",
           855 => x"c9398c08",
           856 => x"fc050880",
           857 => x"2e80c938",
           858 => x"8c088c05",
           859 => x"088c0888",
           860 => x"050826a1",
           861 => x"388c0888",
           862 => x"05088c08",
           863 => x"8c050831",
           864 => x"8c088805",
           865 => x"0c8c08f8",
           866 => x"05088c08",
           867 => x"fc050807",
           868 => x"8c08f805",
           869 => x"0c8c08fc",
           870 => x"0508812a",
           871 => x"8c08fc05",
           872 => x"0c8c088c",
           873 => x"0508812a",
           874 => x"8c088c05",
           875 => x"0cffaf39",
           876 => x"8c089005",
           877 => x"08802e8f",
           878 => x"388c0888",
           879 => x"0508708c",
           880 => x"08f4050c",
           881 => x"518d398c",
           882 => x"08f80508",
           883 => x"708c08f4",
           884 => x"050c518c",
           885 => x"08f40508",
           886 => x"800c853d",
           887 => x"0d8c0c04",
           888 => x"fd3d0d80",
           889 => x"0b9e9808",
           890 => x"54547281",
           891 => x"2e983873",
           892 => x"a6fc0ced",
           893 => x"aa3fec88",
           894 => x"3f9fac52",
           895 => x"8151eee1",
           896 => x"3f800851",
           897 => x"9e3f72a6",
           898 => x"fc0ced93",
           899 => x"3febf13f",
           900 => x"9fac5281",
           901 => x"51eeca3f",
           902 => x"80085187",
           903 => x"3f00ff39",
           904 => x"00ff39f7",
           905 => x"3d0d7b9f",
           906 => x"b00882c8",
           907 => x"11085a54",
           908 => x"5a77802e",
           909 => x"80d93881",
           910 => x"88188419",
           911 => x"08ff0581",
           912 => x"712b5955",
           913 => x"59807424",
           914 => x"80e93880",
           915 => x"7424b538",
           916 => x"73822b78",
           917 => x"11880556",
           918 => x"56818019",
           919 => x"08770653",
           920 => x"72802eb5",
           921 => x"38781670",
           922 => x"08535379",
           923 => x"51740853",
           924 => x"722dff14",
           925 => x"fc17fc17",
           926 => x"79812c5a",
           927 => x"57575473",
           928 => x"8025d638",
           929 => x"77085877",
           930 => x"ffad389f",
           931 => x"b00853bc",
           932 => x"1308a538",
           933 => x"7951ff85",
           934 => x"3f740853",
           935 => x"722dff14",
           936 => x"fc17fc17",
           937 => x"79812c5a",
           938 => x"57575473",
           939 => x"8025ffa9",
           940 => x"38d23980",
           941 => x"57ff9439",
           942 => x"7251bc13",
           943 => x"0853722d",
           944 => x"7951fed9",
           945 => x"3fff3d0d",
           946 => x"a6b40bfc",
           947 => x"05700852",
           948 => x"5270ff2e",
           949 => x"9138702d",
           950 => x"fc127008",
           951 => x"525270ff",
           952 => x"2e098106",
           953 => x"f138833d",
           954 => x"0d0404ec",
           955 => x"943f0400",
           956 => x"00ffffff",
           957 => x"ff00ffff",
           958 => x"ffff00ff",
           959 => x"ffffff00",
           960 => x"00000040",
           961 => x"64756d6d",
           962 => x"792e6578",
           963 => x"65000000",
           964 => x"43000000",
           965 => x"00000000",
           966 => x"00000000",
           967 => x"00000000",
           968 => x"0000133c",
           969 => x"00008004",
           970 => x"00008008",
           971 => x"0000800c",
           972 => x"00008010",
           973 => x"00008014",
           974 => x"00008018",
           975 => x"0000801c",
           976 => x"00008020",
           977 => x"00008030",
           978 => x"0000a004",
           979 => x"0000a008",
           980 => x"0000a00c",
           981 => x"0000a010",
           982 => x"0000a014",
           983 => x"0000a020",
           984 => x"0000a024",
           985 => x"0000a028",
           986 => x"0000a02c",
           987 => x"0000a030",
           988 => x"0000a034",
           989 => x"0000a038",
           990 => x"0000a03c",
           991 => x"0000e004",
           992 => x"0000e008",
           993 => x"0000e00c",
           994 => x"0000e010",
           995 => x"00000000",
           996 => x"00000000",
           997 => x"00000000",
           998 => x"00000000",
           999 => x"00000000",
          1000 => x"00000000",
          1001 => x"00000000",
          1002 => x"00000000",
          1003 => x"00000f04",
          1004 => x"00000fb4",
          1005 => x"00000000",
          1006 => x"0000121c",
          1007 => x"00001278",
          1008 => x"000012d4",
          1009 => x"00000000",
          1010 => x"00000000",
          1011 => x"00000000",
          1012 => x"00000000",
          1013 => x"00000000",
          1014 => x"00000000",
          1015 => x"00000000",
          1016 => x"00000000",
          1017 => x"00000000",
          1018 => x"00000f10",
          1019 => x"00000000",
          1020 => x"00000000",
          1021 => x"00000000",
          1022 => x"00000000",
          1023 => x"00000000",
          1024 => x"00000000",
          1025 => x"00000000",
          1026 => x"00000000",
          1027 => x"00000000",
          1028 => x"00000000",
          1029 => x"00000000",
          1030 => x"00000000",
          1031 => x"00000000",
          1032 => x"00000000",
          1033 => x"00000000",
          1034 => x"00000000",
          1035 => x"00000000",
          1036 => x"00000000",
          1037 => x"00000000",
          1038 => x"00000000",
          1039 => x"00000000",
          1040 => x"00000000",
          1041 => x"00000000",
          1042 => x"00000000",
          1043 => x"00000000",
          1044 => x"00000000",
          1045 => x"00000000",
          1046 => x"00000000",
          1047 => x"00000001",
          1048 => x"330eabcd",
          1049 => x"1234e66d",
          1050 => x"deec0005",
          1051 => x"000b0000",
          1052 => x"00000000",
          1053 => x"00000000",
          1054 => x"00000000",
          1055 => x"00000000",
          1056 => x"00000000",
          1057 => x"00000000",
          1058 => x"00000000",
          1059 => x"00000000",
          1060 => x"00000000",
          1061 => x"00000000",
          1062 => x"00000000",
          1063 => x"00000000",
          1064 => x"00000000",
          1065 => x"00000000",
          1066 => x"00000000",
          1067 => x"00000000",
          1068 => x"00000000",
          1069 => x"00000000",
          1070 => x"00000000",
          1071 => x"00000000",
          1072 => x"00000000",
          1073 => x"00000000",
          1074 => x"00000000",
          1075 => x"00000000",
          1076 => x"00000000",
          1077 => x"00000000",
          1078 => x"00000000",
          1079 => x"00000000",
          1080 => x"00000000",
          1081 => x"00000000",
          1082 => x"00000000",
          1083 => x"00000000",
          1084 => x"00000000",
          1085 => x"00000000",
          1086 => x"00000000",
          1087 => x"00000000",
          1088 => x"00000000",
          1089 => x"00000000",
          1090 => x"00000000",
          1091 => x"00000000",
          1092 => x"00000000",
          1093 => x"00000000",
          1094 => x"00000000",
          1095 => x"00000000",
          1096 => x"00000000",
          1097 => x"00000000",
          1098 => x"00000000",
          1099 => x"00000000",
          1100 => x"00000000",
          1101 => x"00000000",
          1102 => x"00000000",
          1103 => x"00000000",
          1104 => x"00000000",
          1105 => x"00000000",
          1106 => x"00000000",
          1107 => x"00000000",
          1108 => x"00000000",
          1109 => x"00000000",
          1110 => x"00000000",
          1111 => x"00000000",
          1112 => x"00000000",
          1113 => x"00000000",
          1114 => x"00000000",
          1115 => x"00000000",
          1116 => x"00000000",
          1117 => x"00000000",
          1118 => x"00000000",
          1119 => x"00000000",
          1120 => x"00000000",
          1121 => x"00000000",
          1122 => x"00000000",
          1123 => x"00000000",
          1124 => x"00000000",
          1125 => x"00000000",
          1126 => x"00000000",
          1127 => x"00000000",
          1128 => x"00000000",
          1129 => x"00000000",
          1130 => x"00000000",
          1131 => x"00000000",
          1132 => x"00000000",
          1133 => x"00000000",
          1134 => x"00000000",
          1135 => x"00000000",
          1136 => x"00000000",
          1137 => x"00000000",
          1138 => x"00000000",
          1139 => x"00000000",
          1140 => x"00000000",
          1141 => x"00000000",
          1142 => x"00000000",
          1143 => x"00000000",
          1144 => x"00000000",
          1145 => x"00000000",
          1146 => x"00000000",
          1147 => x"00000000",
          1148 => x"00000000",
          1149 => x"00000000",
          1150 => x"00000000",
          1151 => x"00000000",
          1152 => x"00000000",
          1153 => x"00000000",
          1154 => x"00000000",
          1155 => x"00000000",
          1156 => x"00000000",
          1157 => x"00000000",
          1158 => x"00000000",
          1159 => x"00000000",
          1160 => x"00000000",
          1161 => x"00000000",
          1162 => x"00000000",
          1163 => x"00000000",
          1164 => x"00000000",
          1165 => x"00000000",
          1166 => x"00000000",
          1167 => x"00000000",
          1168 => x"00000000",
          1169 => x"00000000",
          1170 => x"00000000",
          1171 => x"00000000",
          1172 => x"00000000",
          1173 => x"00000000",
          1174 => x"00000000",
          1175 => x"00000000",
          1176 => x"00000000",
          1177 => x"00000000",
          1178 => x"00000000",
          1179 => x"00000000",
          1180 => x"00000000",
          1181 => x"00000000",
          1182 => x"00000000",
          1183 => x"00000000",
          1184 => x"00000000",
          1185 => x"00000000",
          1186 => x"00000000",
          1187 => x"00000000",
          1188 => x"00000000",
          1189 => x"00000000",
          1190 => x"00000000",
          1191 => x"00000000",
          1192 => x"00000000",
          1193 => x"00000000",
          1194 => x"00000000",
          1195 => x"00000000",
          1196 => x"00000000",
          1197 => x"00000000",
          1198 => x"00000000",
          1199 => x"00000000",
          1200 => x"00000000",
          1201 => x"00000000",
          1202 => x"00000000",
          1203 => x"00000000",
          1204 => x"00000000",
          1205 => x"00000000",
          1206 => x"00000000",
          1207 => x"00000000",
          1208 => x"00000000",
          1209 => x"00000000",
          1210 => x"00000000",
          1211 => x"00000000",
          1212 => x"00000000",
          1213 => x"00000000",
          1214 => x"00000000",
          1215 => x"00000000",
          1216 => x"00000000",
          1217 => x"00000000",
          1218 => x"00000000",
          1219 => x"00000000",
          1220 => x"00000000",
          1221 => x"00000000",
          1222 => x"00000000",
          1223 => x"00000000",
          1224 => x"00000000",
          1225 => x"00000000",
          1226 => x"00000000",
          1227 => x"00000000",
          1228 => x"ffffffff",
          1229 => x"00000000",
          1230 => x"ffffffff",
          1231 => x"00000000",
          1232 => x"00000000",

        others => x"00000000"
    );

begin
    process (clk) begin
        if (clk'event and clk = '1') then
            if (memAWriteEnable = '1') and (memBWriteEnable = '1') and (memAAddr=memBAddr) and (memAWrite/=memBWrite) then
                report "write collision" severity failure;
            end if;

            if (memAWriteEnable = '1') then
                ram(to_integer(unsigned(memAAddr))) := memAWrite;
                memARead <= memAWrite;
            else
                memARead <= ram(to_integer(unsigned(memAAddr)));
            end if;
        end if;
    end process;

    process (clk) begin
        if (clk'event and clk = '1') then
            if (memBWriteEnable = '1') then
                ram(to_integer(unsigned(memBAddr))) := memBWrite;
                memBRead <= memBWrite;
            else
                memBRead <= ram(to_integer(unsigned(memBAddr)));
            end if;
        end if;
    end process;



end dualport_ram_arch;